VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO mp_cache_data_array
   CLASS BLOCK ;
   SIZE 893.29 BY 106.0125 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
      END
   END din0[199]
   PIN din0[200]
      DIRECTION INPUT ;
      PORT
      END
   END din0[200]
   PIN din0[201]
      DIRECTION INPUT ;
      PORT
      END
   END din0[201]
   PIN din0[202]
      DIRECTION INPUT ;
      PORT
      END
   END din0[202]
   PIN din0[203]
      DIRECTION INPUT ;
      PORT
      END
   END din0[203]
   PIN din0[204]
      DIRECTION INPUT ;
      PORT
      END
   END din0[204]
   PIN din0[205]
      DIRECTION INPUT ;
      PORT
      END
   END din0[205]
   PIN din0[206]
      DIRECTION INPUT ;
      PORT
      END
   END din0[206]
   PIN din0[207]
      DIRECTION INPUT ;
      PORT
      END
   END din0[207]
   PIN din0[208]
      DIRECTION INPUT ;
      PORT
      END
   END din0[208]
   PIN din0[209]
      DIRECTION INPUT ;
      PORT
      END
   END din0[209]
   PIN din0[210]
      DIRECTION INPUT ;
      PORT
      END
   END din0[210]
   PIN din0[211]
      DIRECTION INPUT ;
      PORT
      END
   END din0[211]
   PIN din0[212]
      DIRECTION INPUT ;
      PORT
      END
   END din0[212]
   PIN din0[213]
      DIRECTION INPUT ;
      PORT
      END
   END din0[213]
   PIN din0[214]
      DIRECTION INPUT ;
      PORT
      END
   END din0[214]
   PIN din0[215]
      DIRECTION INPUT ;
      PORT
      END
   END din0[215]
   PIN din0[216]
      DIRECTION INPUT ;
      PORT
      END
   END din0[216]
   PIN din0[217]
      DIRECTION INPUT ;
      PORT
      END
   END din0[217]
   PIN din0[218]
      DIRECTION INPUT ;
      PORT
      END
   END din0[218]
   PIN din0[219]
      DIRECTION INPUT ;
      PORT
      END
   END din0[219]
   PIN din0[220]
      DIRECTION INPUT ;
      PORT
      END
   END din0[220]
   PIN din0[221]
      DIRECTION INPUT ;
      PORT
      END
   END din0[221]
   PIN din0[222]
      DIRECTION INPUT ;
      PORT
      END
   END din0[222]
   PIN din0[223]
      DIRECTION INPUT ;
      PORT
      END
   END din0[223]
   PIN din0[224]
      DIRECTION INPUT ;
      PORT
      END
   END din0[224]
   PIN din0[225]
      DIRECTION INPUT ;
      PORT
      END
   END din0[225]
   PIN din0[226]
      DIRECTION INPUT ;
      PORT
      END
   END din0[226]
   PIN din0[227]
      DIRECTION INPUT ;
      PORT
      END
   END din0[227]
   PIN din0[228]
      DIRECTION INPUT ;
      PORT
      END
   END din0[228]
   PIN din0[229]
      DIRECTION INPUT ;
      PORT
      END
   END din0[229]
   PIN din0[230]
      DIRECTION INPUT ;
      PORT
      END
   END din0[230]
   PIN din0[231]
      DIRECTION INPUT ;
      PORT
      END
   END din0[231]
   PIN din0[232]
      DIRECTION INPUT ;
      PORT
      END
   END din0[232]
   PIN din0[233]
      DIRECTION INPUT ;
      PORT
      END
   END din0[233]
   PIN din0[234]
      DIRECTION INPUT ;
      PORT
      END
   END din0[234]
   PIN din0[235]
      DIRECTION INPUT ;
      PORT
      END
   END din0[235]
   PIN din0[236]
      DIRECTION INPUT ;
      PORT
      END
   END din0[236]
   PIN din0[237]
      DIRECTION INPUT ;
      PORT
      END
   END din0[237]
   PIN din0[238]
      DIRECTION INPUT ;
      PORT
      END
   END din0[238]
   PIN din0[239]
      DIRECTION INPUT ;
      PORT
      END
   END din0[239]
   PIN din0[240]
      DIRECTION INPUT ;
      PORT
      END
   END din0[240]
   PIN din0[241]
      DIRECTION INPUT ;
      PORT
      END
   END din0[241]
   PIN din0[242]
      DIRECTION INPUT ;
      PORT
      END
   END din0[242]
   PIN din0[243]
      DIRECTION INPUT ;
      PORT
      END
   END din0[243]
   PIN din0[244]
      DIRECTION INPUT ;
      PORT
      END
   END din0[244]
   PIN din0[245]
      DIRECTION INPUT ;
      PORT
      END
   END din0[245]
   PIN din0[246]
      DIRECTION INPUT ;
      PORT
      END
   END din0[246]
   PIN din0[247]
      DIRECTION INPUT ;
      PORT
      END
   END din0[247]
   PIN din0[248]
      DIRECTION INPUT ;
      PORT
      END
   END din0[248]
   PIN din0[249]
      DIRECTION INPUT ;
      PORT
      END
   END din0[249]
   PIN din0[250]
      DIRECTION INPUT ;
      PORT
      END
   END din0[250]
   PIN din0[251]
      DIRECTION INPUT ;
      PORT
      END
   END din0[251]
   PIN din0[252]
      DIRECTION INPUT ;
      PORT
      END
   END din0[252]
   PIN din0[253]
      DIRECTION INPUT ;
      PORT
      END
   END din0[253]
   PIN din0[254]
      DIRECTION INPUT ;
      PORT
      END
   END din0[254]
   PIN din0[255]
      DIRECTION INPUT ;
      PORT
      END
   END din0[255]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[7]
   PIN wmask0[8]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[8]
   PIN wmask0[9]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[9]
   PIN wmask0[10]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[10]
   PIN wmask0[11]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[11]
   PIN wmask0[12]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[12]
   PIN wmask0[13]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[13]
   PIN wmask0[14]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[14]
   PIN wmask0[15]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[15]
   PIN wmask0[16]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[16]
   PIN wmask0[17]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[17]
   PIN wmask0[18]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[18]
   PIN wmask0[19]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[19]
   PIN wmask0[20]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[20]
   PIN wmask0[21]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[21]
   PIN wmask0[22]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[22]
   PIN wmask0[23]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[23]
   PIN wmask0[24]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[24]
   PIN wmask0[25]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[25]
   PIN wmask0[26]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[26]
   PIN wmask0[27]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[27]
   PIN wmask0[28]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[28]
   PIN wmask0[29]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[29]
   PIN wmask0[30]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[30]
   PIN wmask0[31]
      DIRECTION INPUT ;
      PORT
      END
   END wmask0[31]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[79]
   PIN dout0[80]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[80]
   PIN dout0[81]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[81]
   PIN dout0[82]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[82]
   PIN dout0[83]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[83]
   PIN dout0[84]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[84]
   PIN dout0[85]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[85]
   PIN dout0[86]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[86]
   PIN dout0[87]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[87]
   PIN dout0[88]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[88]
   PIN dout0[89]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[89]
   PIN dout0[90]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[90]
   PIN dout0[91]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[91]
   PIN dout0[92]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[92]
   PIN dout0[93]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[93]
   PIN dout0[94]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[94]
   PIN dout0[95]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[95]
   PIN dout0[96]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[96]
   PIN dout0[97]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[97]
   PIN dout0[98]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[98]
   PIN dout0[99]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[99]
   PIN dout0[100]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[100]
   PIN dout0[101]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[101]
   PIN dout0[102]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[102]
   PIN dout0[103]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[103]
   PIN dout0[104]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[104]
   PIN dout0[105]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[105]
   PIN dout0[106]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[106]
   PIN dout0[107]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[107]
   PIN dout0[108]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[108]
   PIN dout0[109]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[109]
   PIN dout0[110]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[110]
   PIN dout0[111]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[111]
   PIN dout0[112]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[112]
   PIN dout0[113]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[113]
   PIN dout0[114]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[114]
   PIN dout0[115]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[115]
   PIN dout0[116]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[116]
   PIN dout0[117]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[117]
   PIN dout0[118]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[118]
   PIN dout0[119]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[119]
   PIN dout0[120]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[120]
   PIN dout0[121]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[121]
   PIN dout0[122]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[122]
   PIN dout0[123]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[123]
   PIN dout0[124]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[124]
   PIN dout0[125]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[125]
   PIN dout0[126]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[126]
   PIN dout0[127]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[127]
   PIN dout0[128]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[128]
   PIN dout0[129]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[129]
   PIN dout0[130]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[130]
   PIN dout0[131]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[131]
   PIN dout0[132]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[132]
   PIN dout0[133]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[133]
   PIN dout0[134]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[134]
   PIN dout0[135]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[135]
   PIN dout0[136]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[136]
   PIN dout0[137]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[137]
   PIN dout0[138]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[138]
   PIN dout0[139]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[139]
   PIN dout0[140]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[140]
   PIN dout0[141]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[141]
   PIN dout0[142]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[142]
   PIN dout0[143]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[143]
   PIN dout0[144]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[144]
   PIN dout0[145]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[145]
   PIN dout0[146]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[146]
   PIN dout0[147]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[147]
   PIN dout0[148]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[148]
   PIN dout0[149]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[149]
   PIN dout0[150]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[150]
   PIN dout0[151]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[151]
   PIN dout0[152]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[152]
   PIN dout0[153]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[153]
   PIN dout0[154]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[154]
   PIN dout0[155]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[155]
   PIN dout0[156]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[156]
   PIN dout0[157]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[157]
   PIN dout0[158]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[158]
   PIN dout0[159]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[159]
   PIN dout0[160]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[160]
   PIN dout0[161]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[161]
   PIN dout0[162]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[162]
   PIN dout0[163]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[163]
   PIN dout0[164]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[164]
   PIN dout0[165]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[165]
   PIN dout0[166]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[166]
   PIN dout0[167]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[167]
   PIN dout0[168]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[168]
   PIN dout0[169]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[169]
   PIN dout0[170]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[170]
   PIN dout0[171]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[171]
   PIN dout0[172]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[172]
   PIN dout0[173]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[173]
   PIN dout0[174]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[174]
   PIN dout0[175]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[175]
   PIN dout0[176]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[176]
   PIN dout0[177]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[177]
   PIN dout0[178]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[178]
   PIN dout0[179]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[179]
   PIN dout0[180]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[180]
   PIN dout0[181]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[181]
   PIN dout0[182]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[182]
   PIN dout0[183]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[183]
   PIN dout0[184]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[184]
   PIN dout0[185]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[185]
   PIN dout0[186]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[186]
   PIN dout0[187]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[187]
   PIN dout0[188]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[188]
   PIN dout0[189]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[189]
   PIN dout0[190]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[190]
   PIN dout0[191]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[191]
   PIN dout0[192]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[192]
   PIN dout0[193]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[193]
   PIN dout0[194]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[194]
   PIN dout0[195]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[195]
   PIN dout0[196]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[196]
   PIN dout0[197]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[197]
   PIN dout0[198]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[198]
   PIN dout0[199]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[199]
   PIN dout0[200]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[200]
   PIN dout0[201]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[201]
   PIN dout0[202]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[202]
   PIN dout0[203]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[203]
   PIN dout0[204]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[204]
   PIN dout0[205]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[205]
   PIN dout0[206]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[206]
   PIN dout0[207]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[207]
   PIN dout0[208]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[208]
   PIN dout0[209]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[209]
   PIN dout0[210]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[210]
   PIN dout0[211]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[211]
   PIN dout0[212]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[212]
   PIN dout0[213]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[213]
   PIN dout0[214]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[214]
   PIN dout0[215]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[215]
   PIN dout0[216]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[216]
   PIN dout0[217]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[217]
   PIN dout0[218]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[218]
   PIN dout0[219]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[219]
   PIN dout0[220]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[220]
   PIN dout0[221]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[221]
   PIN dout0[222]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[222]
   PIN dout0[223]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[223]
   PIN dout0[224]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[224]
   PIN dout0[225]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[225]
   PIN dout0[226]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[226]
   PIN dout0[227]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[227]
   PIN dout0[228]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[228]
   PIN dout0[229]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[229]
   PIN dout0[230]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[230]
   PIN dout0[231]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[231]
   PIN dout0[232]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[232]
   PIN dout0[233]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[233]
   PIN dout0[234]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[234]
   PIN dout0[235]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[235]
   PIN dout0[236]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[236]
   PIN dout0[237]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[237]
   PIN dout0[238]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[238]
   PIN dout0[239]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[239]
   PIN dout0[240]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[240]
   PIN dout0[241]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[241]
   PIN dout0[242]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[242]
   PIN dout0[243]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[243]
   PIN dout0[244]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[244]
   PIN dout0[245]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[245]
   PIN dout0[246]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[246]
   PIN dout0[247]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[247]
   PIN dout0[248]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[248]
   PIN dout0[249]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[249]
   PIN dout0[250]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[250]
   PIN dout0[251]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[251]
   PIN dout0[252]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[252]
   PIN dout0[253]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[253]
   PIN dout0[254]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[254]
   PIN dout0[255]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[255]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 893.15 105.8725 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 893.15 105.8725 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 893.15 105.8725 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 893.15 105.8725 ;
   END
END    mp_cache_data_array
END    LIBRARY
