VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO mp_cache_tag_array
   CLASS BLOCK ;
   SIZE 84.515 BY 46.5 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
      END
   END din0[22]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
      END
   END dout0[22]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 84.375 46.36 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 84.375 46.36 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 84.375 46.36 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 84.375 46.36 ;
   END
END    mp_cache_tag_array
END    LIBRARY
